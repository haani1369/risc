`default_nettype none


module reorder_buffer (
  input wire clk_in,
  input wire rst_in,

  
);



endmodule


`default_nettype wire
