`default_nettype none

module writeback (

);

endmodule

`default_nettype wire
